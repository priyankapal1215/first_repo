module tb;
initial begin
	$display("hello world");
end
endmodule
